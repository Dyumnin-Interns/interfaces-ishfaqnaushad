module dut(CLK,
	   RST_N,

	   write_address,
	   write_data,
	   write_en,
	   write_rdy,

	   read_address,
	   read_en,
	   read_data,
	   read_rdy);
  dut test(
